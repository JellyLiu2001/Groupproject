Untitled Sketch
R8 0 11 220
S2 8 83 control_S2 0 generic_switch OFF
VS2 control_S2 0 DC 0
R3 0 8 220
R2 0 8 220
R7 16 13 220
R1 0 8 220
R4 0 8 220
S5_1 17 8 control_S5_1 0 generic_switch OFF
S5_2 11 8 control_S5_2 0 generic_switch ON
VS5_1 control_S5_1 0 DC 0
VS5_2 control_S5_2 0 DC 5
R5 12 14 220
S3 8 82 control_S3 0 generic_switch OFF
VS3 control_S3 0 DC 0
S1 8 84 control_S1 0 generic_switch OFF
VS1 control_S1 0 DC 0
R6 15 10 220
S4 8 81 control_S4 0 generic_switch OFF
VS4 control_S4 0 DC 0

.MODEL generic_switch SW(Ron=1m Roff=1Meg Vt=2.5)

.options savecurrents
.OP
*.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END